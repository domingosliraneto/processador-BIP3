LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PC IS
	PORT(E : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 clk, EN, rst : IN STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(10 DOWNTO 0));
END PC;

ARCHITECTURE arch OF PC IS
BEGIN
	PROCESS(E, clk, EN, rst)
	BEGIN
		IF(rst = '1') THEN
			S <= (OTHERS => '0');
		ELSIF(RISING_EDGE(clk)) THEN
			IF(EN = '1') THEN
				S <= E;
			END IF;
		END IF;
	END PROCESS;
END;