LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux2_1 IS
	PORT(E1, E0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  SEL : IN STD_LOGIC;
		  S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END mux2_1;

ARCHITECTURE arch OF mux2_1 IS
BEGIN
	S <= E0 WHEN SEL = '0' ELSE
	     E1;
END;